stabilnosc

vwe 1 0 ac 1
e1 2 0 laplace {v(1)}={ku0/((1+s/1.58k)*(1+s/15.8k)*(1+s/158k))}
.param ku0=100k
.step dec param ku0 10 10k 12
.ac dec 10 1 100g
.probe
.end

; Podobniez
; 1. Symulacja
; 2. Performance Analysis -> wizard
; 3. Phase Margin
; 4. phase trace p(v(2))
; 5. magnitude trace in db vdb(2)
; 6. cursor -> sea forw lev -45

; Wynik: ok. 2.2875k