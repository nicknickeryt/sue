zabezpieczenie termicnze

; Zalozenie - temp. pokojowa 20C

.model BC107 NPN(Is=40.72f Bf=407 Vaf=21.03 Ikf=1 Ise=40.72f Ne=1.305 Ikr=3.726
+ Isc=594.8p Nc=2.033 Rc=1.393 Cje=12.5p Vje=.5391 Mje=.4869 Tf=441.1p Cjc=6p
+ Mjc=.3821 Tr=114n Xtb=1.5 )

.model BC547B NPN(IS=2.39E-14 NF=1.008 ISE=3.545E-15 NE=1.541 BF=294.3 IKF=0.1357 
+ VAF=63.2 NR=1.004 ISC=6.272E-14 NC=1.243 BR=7.946 IKR=0.1144 VAR=25.9 RB=1 IRB=1.00E-06 
+ RBM=1 RE=0.4683 RC=0.85 XTB=0 EG=1.11 XTI=3 CJE=1.358E-11 VJE=0.65 MJE=0.3279 TF=4.391E-10 
+ XTF=120 VTF=2.643 ITF=0.7495 PTF=0 CJC=3.728E-12 VJC=0.3997 MJC=0.2955 XCJC=0.6193 TR=1.00E-32 
+ CJS=0 VJS=0.75 MJS=0.333 FC=0.9579)

.model BZX84C12L D(Is=.6n Rs=.5 Cjo=150p nbv=5 bv=12 Ibv=1m)

V vcc 0 30

Q1 vcc 1 out  BC107 
Q2 1 2 0 BC107

D 0 1 BZX84C12L


R1 out 0 1k
R2 2 3 1k
R3 vcc 2 82k
R4 vcc 1 2.2k

.param opornik = 400

R5 3 0 {opornik}


.dc param opornik 400 4700 1;
.probe


; R5  = 20 * temperatura
; temperatura = R5/20
; 90% wartosci nominalnej

; 1. Obliczenie wartosci nominalnej
; R4 = 20 * 20 = 400
; wtedy Vout = 11.607
; 90% to 10.4463
; Szukane R5 = 1016Ohm
; Temperatura = 1016/20 = 50.8

; Zapami�ta�
; Param, przekszta�cenia, temp. pokojowa to 20C
; Szybko liczyc :))