stabilność

vwe 1 0 ac 1
e1 2 0 laplace {v(1)}={26/((1+s/1.58)*(1+s/15.8k)*(1+s/158k))}
.ac dec 10 1 100g
.probe
.end

; Pamieciowka
; 1. Symulacja
; 2. Trace->Eval. Measurement
; 3. GainMargin(p(v(2)), vdb(2))) ok. 72.53
; 4. PhaseMargin(vdb(2), p(v(2))) ok. 92.05